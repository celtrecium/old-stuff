Z   -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    `     `     `                                                                                                                                                                                                                `     `     `     `     `                          `     `     `     `     `                                 `     `     `     `     `                   `                                        `                                                      `                                        `                          `     `     `     `     `                          `                                        `                                                                                                                                                                                           `                                                      `                                        `                   `                                                      `                                 `     `                                                      `     `                          `     `                   `                                        `                   `                                 `     `                                                                                                                                                                                           `                                                      `                                        `                   `                                                      `                          `            `                                                      `            `            `            `                   `                                        `                   `                          `            `                                                                                                                                                                                           `                                                      `     `     `     `     `     `     `                   `                                                      `                   `                   `                                                      `                   `                   `                   `                                        `                   `                   `                   `                                                                                                                                                                                           `                                                      `                                        `                   `                                                      `            `                          `                                                      `                                        `                   `                                        `                   `            `                          `                                                                                                                                                                                           `                                                      `                                        `                   `                                                      `     `                                 `                                                      `                                        `                   `                                        `                   `     `                                 `                                                                                                                                                                                                  `     `     `     `     `                   `                                        `                          `     `     `     `     `                   `                                        `                                                      `                                        `                          `     `     `     `     `                          `                                        `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           `     `                                                                                                                                                                                                                                                   `     `     `     `     `     `                          `     `     `     `     `                                        `     `     `     `                          `     `     `     `     `     `                   `     `     `     `     `     `                   `                                               `                   `                                 `                                                                                                                                                                                                                                                   `     `                                 `                                        `                          `                          `                   `                                                                           `     `                                 `                                               `                   `                          `     `                                                                                                                                                                                                                                                   `     `                                 `                                        `                          `                          `                   `                                                                           `     `                                 `     `     `     `     `                   `                   `                   `            `                                                                                                                                                                                                                                                   `     `                                 `                                        `                          `                          `                   `                                                                           `     `                                 `                                 `            `                   `            `                   `                                                                                                                                                                                                                                                   `     `                                 `                                        `                          `                          `                   `                                                                           `     `                                 `                                 `            `                   `     `                          `                                                                                                                                                                                                                                                   `     `                                        `     `     `     `     `                          `                                 `                          `     `     `     `     `     `                                 `     `                                 `     `     `     `     `                   `                   `                                 `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   `     `     `     `     `     `     `     `                                        `     `     `                                               `     `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                              `     `     `                                               `     `                                        `     `                                        `     `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                              `     `                                                                                                              `     `                                 `     `     `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                              `     `                                                                                                              `     `                          `     `            `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                              `     `                                                                                                              `     `                   `     `                   `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                              `     `                                                                                                              `     `            `     `                          `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                              `     `                                                                                                              `     `     `     `                                 `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                                     `     `     `                                               `     `                                        `     `     `                                        `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   `     `     `     `     `     `     `     `                                        `     `     `                                               `     `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  