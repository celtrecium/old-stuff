2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         `    `    `    `    `                                                                                                                                                                                                                                                                                                                        `                  `                  `                                                                                                                                                                                                                                                                                                                 `                  `                  `                                                                                                                                                                                                                                                                                                                 `                  `                  `                  `                  `                  `           `                         `    `                                                                                                                                                                                                        `    `    `    `    `                         `                  `                  `    `                         `                                                                                                                                                                                                                                    `                                              `    `    `                  `           `                         `    `                                                                                                                                                                                                                                                                                     `                                                                                                                                                                                                                                                                                                                                                           `                                                                                                                                                                                                                                                                                                                                             `    `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  